module dumpfile;
    initial
    begin
        // $dumpfile("test.vcd");
        // $dumpvars(0,ram_512_tb);
    end
endmodule