`timescale 1 ns/10 ps

module or_16_tb;
    reg [15:0] in_a, in_b, out;
    reg [15:0] rand_in_a, rand_in_b, expected_out;
    localparam period = 20;
    or_16 UUT (.in_a(in_a), .in_b(in_b), .out(out));
    
    initial
    begin
        for (int i = 0; i < 16; i++) begin
            rand_in_a = $urandom();
            rand_in_b = $urandom();
            in_a <= rand_in_a;
            in_b <= rand_in_b;
            #period
            expected_out = rand_in_a | rand_in_b;
            assert(out == expected_out) else begin
                $display("in_a: ", "%b", in_a, ", in_b: ", "%b", in_b, ", out: ", "%b", out, ", expected out: ", "%b", expected_out);
                $fatal(1);
            end;
        end
    end
endmodule
